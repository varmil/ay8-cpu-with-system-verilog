module memory();

endmodule
